module d_ff(d,clk,rst,q);
input d,clk,rst;
output q;
always @(negedge clk or posedge rst)
	



module ripplecounter3();

