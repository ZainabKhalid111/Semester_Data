library verilog;
use verilog.vl_types.all;
entity tst_fsm_lock is
end tst_fsm_lock;
