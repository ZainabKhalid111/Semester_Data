library verilog;
use verilog.vl_types.all;
entity tst_lock is
end tst_lock;
