library verilog;
use verilog.vl_types.all;
entity problem_01 is
end problem_01;
