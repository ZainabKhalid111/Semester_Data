library verilog;
use verilog.vl_types.all;
entity top_johnson is
end top_johnson;
