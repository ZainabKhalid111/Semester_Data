library verilog;
use verilog.vl_types.all;
entity tst_traffic_lights1 is
end tst_traffic_lights1;
