library verilog;
use verilog.vl_types.all;
entity top_for_task_01 is
end top_for_task_01;
