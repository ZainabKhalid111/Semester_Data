library verilog;
use verilog.vl_types.all;
entity test_ripple_adder_4bit is
end test_ripple_adder_4bit;
