library verilog;
use verilog.vl_types.all;
entity test_fa is
end test_fa;
