library verilog;
use verilog.vl_types.all;
entity test_ha2 is
end test_ha2;
