library verilog;
use verilog.vl_types.all;
entity ram_16x8_ex1_testbench is
end ram_16x8_ex1_testbench;
