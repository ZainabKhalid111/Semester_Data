library verilog;
use verilog.vl_types.all;
entity top_level is
end top_level;
