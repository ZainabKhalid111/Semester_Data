library verilog;
use verilog.vl_types.all;
entity tst_fsm_moore is
end tst_fsm_moore;
