library verilog;
use verilog.vl_types.all;
entity stim_fa is
end stim_fa;
