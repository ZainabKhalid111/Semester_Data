library verilog;
use verilog.vl_types.all;
entity top_mux is
end top_mux;
