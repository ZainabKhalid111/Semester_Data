library verilog;
use verilog.vl_types.all;
entity electlocktest is
end electlocktest;
