library verilog;
use verilog.vl_types.all;
entity tst_rom_v2 is
end tst_rom_v2;
