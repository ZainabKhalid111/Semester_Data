library verilog;
use verilog.vl_types.all;
entity test_rippleadder is
end test_rippleadder;
