library verilog;
use verilog.vl_types.all;
entity top_l is
end top_l;
