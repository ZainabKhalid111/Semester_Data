library verilog;
use verilog.vl_types.all;
entity top_counter is
end top_counter;
