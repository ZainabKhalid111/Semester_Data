library verilog;
use verilog.vl_types.all;
entity bcd_top_level is
end bcd_top_level;
