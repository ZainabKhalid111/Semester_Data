library verilog;
use verilog.vl_types.all;
entity tst_rom_32x8 is
end tst_rom_32x8;
