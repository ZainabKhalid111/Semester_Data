library verilog;
use verilog.vl_types.all;
entity stim_rca is
end stim_rca;
