library verilog;
use verilog.vl_types.all;
entity tst_parity_det1 is
end tst_parity_det1;
