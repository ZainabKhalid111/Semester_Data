library verilog;
use verilog.vl_types.all;
entity top_rc is
end top_rc;
