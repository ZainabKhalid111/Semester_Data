library verilog;
use verilog.vl_types.all;
entity test_ha is
end test_ha;
