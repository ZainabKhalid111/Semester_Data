library verilog;
use verilog.vl_types.all;
entity three_bcd_top_level is
end three_bcd_top_level;
