library verilog;
use verilog.vl_types.all;
entity stim_ripple is
end stim_ripple;
