library verilog;
use verilog.vl_types.all;
entity test_fa1 is
end test_fa1;
