library verilog;
use verilog.vl_types.all;
entity tst_rom_16x8 is
end tst_rom_16x8;
