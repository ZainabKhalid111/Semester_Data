library verilog;
use verilog.vl_types.all;
entity test_ha1 is
end test_ha1;
