library verilog;
use verilog.vl_types.all;
entity tst_rom_v1 is
end tst_rom_v1;
